library work;
  context work.cosim_context;
  use work.cosim.all;


entity tb_cosim is
  generic(
    G_SW_GW_FIFO_PATH : string;
    G_GW_SW_FIFO_PATH : string
  );
end entity;


architecture test of tb_cosim is

  signal clk : std_logic := '0';

  signal st : unsigned(71 downto 0) := (others => '1');

  signal req : requester_out_t;
  signal com : completer_out_t;

begin

  clk <= not clk after 0.5 ns;


  cosim_interface(G_SW_GW_FIFO_PATH, G_GW_SW_FIFO_PATH, clk, req, com);


  afbd_main : entity afbd.Main
  port map (
    clk_i => clk,
    rst_i => '0',

    apb_coms_i(0) => req,
    apb_coms_o(0) => com,

    st_i => std_logic_vector(st)
  );


  counters : process (clk) is
  begin
    if rising_edge(clk) then
      st(71 downto 64) <= st(71 downto 64) - 1;
      st(63 downto 32) <= st(63 downto 32) - 1;
    end if;
  end process;

end architecture;
