context cosim_context is
  library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

  library lapb;
    use lapb.apb.all;

  library ltypes;
    use ltypes.types.all;

  library afbd;
    use afbd.apb;
    use afbd.apb.all;

end context;
